module CPU()

RegFile cpu_regs(clock, reset, raA, raB, wa, wen, wd, rdA, rdB);


endmodule